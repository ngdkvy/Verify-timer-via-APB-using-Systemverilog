package test_pkg;

  import timer_pkg::*;

  `include "base_test.sv"
  `include "reg_def_test.sv"
  `include "reg_rw_test.sv"
  `include "reg_rs_test.sv"
  `include "reg_reserved_test.sv"
  `include "reg_tsr_test.sv"
  `include "cnt_up_div1_test.sv"
  `include "cnt_up_div2_test.sv"
  `include "cnt_up_div4_test.sv"
  `include "cnt_up_div8_test.sv"
  `include "cnt_up_rd_div1_test.sv"
  `include "cnt_up_rd_div2_test.sv"
  `include "cnt_up_rd_div4_test.sv"
  `include "cnt_up_rd_div8_test.sv"
  `include "cnt_up_change_test.sv"
  `include "cnt_dw_div1_test.sv"
  `include "cnt_dw_div2_test.sv"
  `include "cnt_dw_div4_test.sv"
  `include "cnt_dw_div8_test.sv"
  `include "cnt_dw_rd_div1_test.sv"
  `include "cnt_dw_rd_div2_test.sv"
  `include "cnt_dw_rd_div4_test.sv"
  `include "cnt_dw_rd_div8_test.sv"
  `include "cnt_dw_change_test.sv"
  `include "cnt_up_dw_test.sv"
  `include "cnt_up_dw_rd_test.sv"
  `include "cnt_dw_up_test.sv"
  `include "cnt_dw_up_rd_test.sv"
  `include "cnt_up_div_1_8_test.sv"
  `include "cnt_up_div_2_8_test.sv"
  `include "cnt_up_div_4_8_test.sv"
  `include "cnt_dw_div_1_8_test.sv"
  `include "cnt_dw_div_2_8_test.sv"
  `include "cnt_dw_div_4_8_test.sv"
  `include "underflow_en_test.sv"
  `include "underflow_dis_test.sv"
  `include "overflow_en_test.sv"
  `include "overflow_dis_test.sv"
  `include "ud_over_en_test.sv"
  `include "ud_over_dis_test.sv"
endpackage
